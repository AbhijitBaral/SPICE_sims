Peak_rectifier (Rectifier with a filter capacitor)

.include ./diode_model.mod

V1    in GND    DC 0 SIN( 0 1 200 0 0 0 0 ) AC 10
D1    in out    DI_1N4007
C1    out GND   100u
*R1    out GND   1k
.end
