.title peak_rectifier
.model __D1 D
+         vj=2
V1 in GND DC 0 SIN( 0 1 1k 0 0 0 ) AC 1  
D1 in out __D1
C1 out GND 10f
.end
