Fixed bias BJT amplifier

.model BC546B npn ( IS=7.59E-15 VAF=73.4 BF=480 IKF=0.0962 NE=1.2665
+ ISE=3.278E-15 IKR=0.03 ISC=2.00E-13 NC=1.2 NR=1 BR=5 RC=0.25 CJC=6.33E-12
+ FC=0.5 MJC=0.33 VJC=0.65 CJE=1.25E-11 MJE=0.55 VJE=0.65 TF=4.26E-10
+ ITF=0.6 VTF=3 XTF=20 RB=100 IRB=0.0001 RBM=10 RE=0.5 TR=1.50E-07)

V2 Vcc GND DC 5
V1 in GND DC 0 SIN( 0 1m 500 0 0 0 ) AC 1  
Cin1 intb in 10u
Cout1 out intc 10u
R3 Vcc intc 10k
R1 Vcc intb 68k
R2 intb GND 10k
Rl1 out GND 100k
Q1 intc intb 0 BC546B

.end
